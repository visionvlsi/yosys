module fa(a,b,cin,sum,co);

input a,b,cin;
output sum,co;

ha ins1(a,b,s1,c1),
   ins2(cin,s1,sum,c2);

orgate ins3(c1,c2,co);


endmodule
